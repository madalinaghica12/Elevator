library IEEE;
use IEEE.STD_LOGIC_1164.all;
use IEEE.STD_LOGIC_ARITH.all;
use IEEE.STD_LOGIC_UNSIGNED.all;

ENTITY INCREMENTARE_DECREMENTARE IS
	PORT( LED : IN STD_LOGIC;
	RESET : IN STD_LOGIC;
	CLK : IN STD_LOGIC;
	
	ETAJ_CURENT : OUT STD_LOGIC_VECTOR(3 DOWNTO 0);
	ETAJ : OUT STD_LOGIC);
END INCREMENTARE_DECREMENTARE;
	
	
	
	
	
	
	
	
	
	
	
	
	
	
	
	
	
	
	
	
	
	
	
	
	
	
	
	
	
	
	
	
	
	
	
	
	
	
	
	
	
	
	