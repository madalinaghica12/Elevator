library IEEE;
use IEEE.STD_LOGIC_1164.all;

ENTITY CAUTARE_ETAJ IS
	PORT( ETAJ_ACTUAL : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
		  CLOCK, RESET : IN STD_LOGIC;
		  INC_PAR_1 : IN STD_LOGIC;
		  INC_PAR_2 : IN STD_LOGIC;
		  CAUTA_MAI_MARE_1 : IN STD_LOGIC;
		  CAUTA_MAI_MARE_2 : IN STD_LOGIC;
		  CAUTA_MAI_MIC_1 : IN STD_LOGIC;
		  CAUTA_MAI_MIC_2 : IN STD_LOGIC;	  
		  ETAJ_MEMORAT : OUT STD_LOGIC_VECTOR(3 DOWNTO 0);
		  SUS : OUT STD_LOGIC;
		  JOS : OUT STD_LOGIC);
END CAUTARE_ETAJ;
	
ARCHITECTURE CAUTARE_ETAJ OF CAUTARE_ETAJ IS

	COMPONENT NUMARATOR_BIDIRECT IS
		PORT( INTR : IN STD_LOGIC_VECTOR( 3 DOWNTO 0);
			  CLOCK : IN STD_LOGIC;  
			  RESET : IN STD_LOGIC;	 
			  INC_PARALELA: IN STD_LOGIC;
			  NUMARA_SUS : IN STD_LOGIC;
			  NUMARA_JOS : IN STD_LOGIC;
			  IESIRE : OUT  STD_LOGIC_VECTOR( 3 DOWNTO 0);
			  SUS : OUT STD_LOGIC;
			  JOS : OUT STD_LOGIC);
	END COMPONENT NUMARATOR_BIDIRECT;
	
	SIGNAL INCARCARE_PARALELA : STD_LOGIC;
	SIGNAL CAUTA_SUS : STD_LOGIC;
	SIGNAL CAUTA_JOS : STD_LOGIC;
	SIGNAL IESIRI : STD_LOGIC_VECTOR(3 DOWNTO 0);	
		
	BEGIN 
		
		INCARCARE_PARALELA <= INC_PAR_1 OR INC_PAR_2;
		CAUTA_SUS <= CAUTA_MAI_MARE_1 OR CAUTA_MAI_MARE_2;
		CAUTA_JOS <= CAUTA_MAI_MIC_1 OR CAUTA_MAI_MIC_2;
		NUM : NUMARATOR_BIDIRECT PORT MAP(ETAJ_ACTUAL, CLOCK, RESET, INCARCARE_PARALELA, CAUTA_SUS, CAUTA_JOS, IESIRI, SUS, JOS);
		ETAJ_MEMORAT <= IESIRI;	 
		
END CAUTARE_ETAJ;