library IEEE;
use IEEE.STD_LOGIC_1164.all; 
use IEEE.STD_LOGIC_UNSIGNED.all;

ENTITY LIFT IS
	PORT( ETAJE : IN  STD_LOGIC_VECTOR(3 DOWNTO 0);
	CLOCK : IN STD_LOGIC;       
	INTERIOR_EXTERIOR : IN STD_LOGIC ;
	SELECTIE_VITEZA : IN STD_LOGIC;
	SENZOR_PERS : IN STD_LOGIC;
	SUS_JOS : IN STD_LOGIC;
	GREUTATE : IN STD_LOGIC;
	INIT : IN STD_LOGIC;   
	USI : IN STD_LOGIC;
	COMANDA : IN STD_LOGIC;
	LED_USI : OUT STD_LOGIC;
	LED_GREUTATE : OUT STD_LOGIC;	 
	ANOZI : OUT STD_LOGIC_VECTOR( 3 DOWNTO 0);
	CATOZI : OUT STD_LOGIC_VECTOR(6 DOWNTO 0)
	);
END LIFT;

ARCHITECTURE LIFT OF LIFT IS   	
	COMPONENT unitatea_de_memorare is
 	 
port (etaje: in std_logic_vector (3 downto 0);

		interior_exterior, sus_jos, clk, stg :in std_logic; 

		comanda: in std_logic;

		etaj_memorat: in std_logic_vector (3 downto 0);

		sus_ext, jos_ext: out std_logic;

		gasit_c: out std_logic);

end COMPONENT unitatea_de_memorare; 	
	
	
	 COMPONENT TIMP IS
		PORT( INCEPUT_TIMP : IN STD_LOGIC;
	      	 CLK : IN STD_LOGIC;     	
		     SFARSIT_TIMP : OUT STD_LOGIC);
	 END COMPONENT TIMP;
	
	
	COMPONENT CAUTARE_ETAJ IS
		PORT( ETAJ_ACTUAL : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
			 CLOCK, RESET : IN STD_LOGIC;
			 INC_PAR_1 : IN STD_LOGIC;
			 INC_PAR_2 : IN STD_LOGIC;
			 CAUTA_MAI_MARE_1 : IN STD_LOGIC;
			 CAUTA_MAI_MARE_2 : IN STD_LOGIC;
			 CAUTA_MAI_MIC_1 : IN STD_LOGIC;
			 CAUTA_MAI_MIC_2 : IN STD_LOGIC;	  
			 ETAJ_MEMORAT : OUT STD_LOGIC_VECTOR(3 DOWNTO 0);
			 SUS : OUT STD_LOGIC;
			 JOS : OUT STD_LOGIC);
	END COMPONENT CAUTARE_ETAJ;	 
		
		
	COMPONENT SENZORI IS
	PORT( SENZOR_PERSOANA : IN STD_LOGIC;
		 SENZOR_GREUTATE : IN STD_LOGIC;    
		 DESCHIS : OUT STD_LOGIC;
		 LED_GREUTATE : OUT STD_LOGIC);   
	END COMPONENT SENZORI;
		
		
	COMPONENT sel_viteza is
	port( V0, V1: IN std_logic;
		F: out std_logic;
		 sl: in std_logic);
	END COMPONENT sel_viteza;	  
		   
		   
	COMPONENT AFISOR IS
	PORT(ETAJ_ACTUAL : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
		CLOCK : IN STD_LOGIC;
		RESET : IN STD_LOGIC;    
		CATOZI_LED :OUT STD_LOGIC_VECTOR (6 DOWNTO 0);	  
		ANOZI : OUT STD_LOGIC_VECTOR (3 DOWNTO 0));   
	END COMPONENT AFISOR;
	
	
	COMPONENT UNITATE_DE_INTARZIERE IS
		PORT( INCEPUT : IN STD_LOGIC;
		 TIMP :IN STD_LOGIC;
		SFARSIT : OUT STD_LOGIC);   
	END COMPONENT UNITATE_DE_INTARZIERE;		 
	
	
	COMPONENT UNITATE_DE_DIRECTIE IS
	PORT( SCHIMBARE_DIRECTIE : IN STD_LOGIC ;
		 CLOCK : IN STD_LOGIC;
		 RESET : IN STD_LOGIC;  
		 DIRECTIE : OUT STD_LOGIC;  
		 N_DIRECTIE : OUT STD_LOGIC); 
	END COMPONENT UNITATE_DE_DIRECTIE; 
	
	
	COMPONENT INCREMENTARE_DECREMENTARE IS
		PORT( LED : IN STD_LOGIC;
		RESET : IN STD_LOGIC;
		CLK : IN STD_LOGIC;
		N_DIRECTIE : IN STD_LOGIC;
		ETAJ_CURENT : OUT STD_LOGIC_VECTOR(3 DOWNTO 0);
		ETAJ : OUT STD_LOGIC); 
	END COMPONENT INCREMENTARE_DECREMENTARE;   
	
	
	COMPONENT UNITATE_DE_DECIZIE IS
		PORT( INTRARE : IN STD_LOGIC_VECTOR(7 downto 0); 
		      CLOCK : IN STD_LOGIC;
			  RESET : IN STD_LOGIC;
			  IESIRE : OUT STD_LOGIC_VECTOR(3 downto 0));
	END COMPONENT UNITATE_DE_DECIZIE;	 
	
	
	COMPONENT Unitate_de_comanda is
		  port(INTRARE : in std_logic_vector(8 downto 0);
		  CLOCK :in std_logic;
		  RESET : in std_logic;
		  IESIRE : out std_logic_vector(8 downto 0));
	end COMPONENT Unitate_de_comanda;   
	
	
	COMPONENT DIVIZOR_DE_FRECVENTA IS
	PORT( CLOCK	: IN STD_LOGIC;
		  RESET : IN STD_LOGIC;  
		  DIVIZOR : OUT STD_LOGIC);     
END COMPONENT DIVIZOR_DE_FRECVENTA;  
	
	
	COMPONENT divizor is
		port( RESET : IN STD_LOGIC;
		      CLOCK : IN STD_LOGIC;
			  DIVIZOR :	OUT STD_LOGIC);               
	END COMPONENT DIVIZOR;	

signal INTRARE : STD_LOGIC_VECTOR (8 DOWNTO 0);
signal DECIZIE_INCEPUT : STD_LOGIC_VECTOR (7 DOWNTO 0);	
signal IESIRE : STD_LOGIC_VECTOR (8 DOWNTO 0);
signal DECIZIE_FINAL : STD_LOGIC_VECTOR (3 DOWNTO 0);
SIGNAL etaj_memorat : STD_LOGIC_VECTOR(3 DOWNTO 0);
SIGNAL ETAJ_CURENT : STD_LOGIC_VECTOR(3 DOWNTO 0);
SIGNAL SUS,JOS,SUS_EXT,JOS_EXT : STD_LOGIC;
SIGNAL COMANDA1, DESCHIS: STD_LOGIC;	 
SIGNAL N_DIRECTIE, DIRECTIE : STD_LOGIC;		   
SIGNAL SFARSIT_TIMP, SFARSIT : STD_LOGIC;
SIGNAL CLK : STD_LOGIC;
SIGNAL INCET, ACCELERAT :STD_LOGIC;	   
SIGNAL ETAJ : STD_LOGIC;


BEGIN
	
	INTRARE(0) <= USI;
	INTRARE(1) <= SFARSIT_TIMP;
	INTRARE(2) <= DESCHIS;		  
	INTRARE(3) <= COMANDA;
	INTRARE(4) <= DIRECTIE;
	INTRARE(5) <= jos; --------
	INTRARE(6) <= sus; ---------
	INTRARE(7) <= DECIZIE_FINAL(0);
	INTRARE(8) <= SFARSIT;		 
	
	
	C1: Unitate_de_comanda PORT MAP(INTRARE,CLOCK,INIT,IESIRE); 
	
	
	DECIZIE_INCEPUT(0) <= IESIRE(2);  ------------
	DECIZIE_INCEPUT(1) <= COMANDA1;	
	DECIZIE_INCEPUT(2) <= DIRECTIE;	  
	DECIZIE_INCEPUT(3) <= SUS_EXT;
	DECIZIE_INCEPUT(4) <= JOS_EXT;
	DECIZIE_INCEPUT(5) <= sus;		-------
	DECIZIE_INCEPUT(6) <= jos;		--------
	DECIZIE_INCEPUT(7) <= ETAJ;	
	
	C2 : UNITATE_DE_DECIZIE port map(DECIZIE_INCEPUT,CLOCK,INIT,DECIZIE_FINAL);
	
	C3 : unitatea_de_memorare PORT MAP(ETAJE,INTERIOR_EXTERIOR,SUS_JOS,CLOCK,IESIRE(0),COMANDA,etaj_memorat, SUS_EXT, JOS_EXT,COMANDA1);
	
	C4 : CAUTARE_ETAJ PORT MAP (ETAJ_CURENT,CLOCK,INIT,IESIRE(6),DECIZIE_FINAL(3),IESIRE(4),DECIZIE_FINAL(1), IESIRE(5), DECIZIE_FINAL(2), ETAJ_MEMORAT,SUS, JOS);
	
	C5 : INCREMENTARE_DECREMENTARE PORT MAP(IESIRE(1),INIT,CLK,N_DIRECTIE,ETAJ_CURENT,ETAJ);
	C6 :  UNITATE_DE_DIRECTIE PORT MAP(IESIRE(3),CLOCK,INIT,DIRECTIE,N_DIRECTIE);
	C7 : TIMP PORT MAP(IESIRE(7),ACCELERAT,SFARSIT_TIMP);
	C8 : SENZORI PORT MAP(SENZOR_PERS,GREUTATE,DESCHIS,LED_GREUTATE);
	C9 : UNITATE_DE_INTARZIERE PORT MAP(IESIRE(8),ACCELERAT,SFARSIT);
	C10 : DIVIZOR_DE_FRECVENTA PORT MAP(CLOCK,INIT,ACCELERAT);
	C11 : divizor  PORT MAP(INIT, CLOCK,INCET) ;
	C12 : SEL_VITEZA PORT MAP  (ACCELERAT,INCET,CLK,SELECTIE_VITEZA);
 	C13 : AFISOR PORT MAP (ETAJ_CURENT,CLOCK,INIT,CATOZI,ANOZI);
	Led_usi	<=	iesire(7);
END LIFT;