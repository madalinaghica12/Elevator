library IEEE;
use IEEE.STD_LOGIC_1164.all;

ENTITY UNITATE_DE_DIRECTIE IS
	PORT( SCHIMBARE_DIRECTIE : IN STD_LOGIC ;
		 CLOCK : IN STD_LOGIC;
		 RESET : IN STD_LOGIC;  
		 DIRECTIE : OUT STD_LOGIC;  
		 N_DIRECTIE : OUT STD_LOGIC); 
END UNITATE_DE_DIRECTIE;

ARCHITECTURE UNITATE_DE_DIRECTIE OF UNITATE_DE_DIRECTIE IS

	COMPONENT BISTABIL_JK IS
		PORT( J : IN STD_LOGIC; 
	   		  K : IN STD_LOGIC; 
		 	 CLOCK : IN STD_LOGIC;   
		 	 Q : OUT STD_LOGIC;
		 	 BQ : OUT STD_LOGIC);  
	END COMPONENT;

	SIGNAL J_DIRECTIE, K_DIRECTIE : STD_LOGIC;
	BEGIN 
		J_DIRECTIE <= SCHIMBARE_DIRECTIE;
		K_DIRECTIE <= SCHIMBARE_DIRECTIE OR RESET;
		BISTABIL : BISTABIL_JK PORT MAP(J_DIRECTIE, K_DIRECTIE, CLOCK, DIRECTIE, N_DIRECTIE); 
		
END UNITATE_DE_DIRECTIE;
	